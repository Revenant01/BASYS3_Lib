`define RESET  3'b000
`define IDLE   3'b001
`define START  3'b011 // transmitter only
`define DATA   3'b010
`define PARITY 3'b110
`define STOP   3'b111